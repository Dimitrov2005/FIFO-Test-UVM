package environment_package;
   import agent_package::*;
`include "Scoreboard.svh"
   