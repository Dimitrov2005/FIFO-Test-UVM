package agnt_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "Transaction.svh"
`include "Sequencer.svh"
`include "Driver.svh"
`include "Monitor.svh"
`include "agent_config.svh"
`include "Agent.svh"
endpackage
   