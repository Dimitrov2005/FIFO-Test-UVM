class DriverR extends uvm_driver();
   