package agent_package;
`include "Driver.svh"
`include "Monitor.svh"
`include "Sequencer.svh"


endpackage // agent_package
   