package env_pkg;
   
import uvm_pkg::*;
import agnt_pkg::*;
`include "uvm_macros.svh"
`include "Scoreboard.svh"
`include "Environment.svh"
`include "environment_config.svh"
   
   
endpackage // environment_package
   
   