package test_pkg;
   
import uvm_pkg::*;
import env_pkg::*;
`include "uvm_macros.svh"
`include "randSeq.svh"
`include "test.svh"
 
   
endpackage